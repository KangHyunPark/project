`timescale 1ns / 1ps

module tb_systolic_input_buffer;
    parameter CLK_PERIOD = 2;
    parameter HALF_CLK_PERIOD = CLK_PERIOD/2;
    
    parameter DATA_WIDTH = 8;
    parameter length = 16;
    
    reg clk;
    reg rstn;
    
    reg [DATA_WIDTH*length-1:0] din;
    wire [DATA_WIDTH*length-1:0] dout;
    
    initial clk = 1'b1;
    always #HALF_CLK_PERIOD clk = ~clk;
    
    initial begin
        rstn = 1'b0;
        
        repeat (100)
        @(posedge clk); 
        
        rstn = 1'b1;   
        
        repeat (100)
        @(posedge clk); 
        
        @(posedge clk) din=128'b00001111000011100000110100001100000010110000101000001001000010000000011100000110000001010000010000000011000000100000000100000000;
        @(posedge clk) din=128'b00011111000111100001110100011100000110110001101000011001000110000001011100010110000101010001010000010011000100100001000100010000;
        @(posedge clk) din=128'b00101111001011100010110100101100001010110010101000101001001010000010011100100110001001010010010000100011001000100010000100100000;
        @(posedge clk) din=128'b00111111001111100011110100111100001110110011101000111001001110000011011100110110001101010011010000110011001100100011000100110000;
        @(posedge clk) din=128'b01001111010011100100110101001100010010110100101001001001010010000100011101000110010001010100010001000011010000100100000101000000;
        @(posedge clk) din=128'b01011111010111100101110101011100010110110101101001011001010110000101011101010110010101010101010001010011010100100101000101010000;
        @(posedge clk) din=128'b01101111011011100110110101101100011010110110101001101001011010000110011101100110011001010110010001100011011000100110000101100000;
        @(posedge clk) din=128'b01111111011111100111110101111100011110110111101001111001011110000111011101110110011101010111010001110011011100100111000101110000;
        @(posedge clk) din=128'b10001111100011101000110110001100100010111000101010001001100010001000011110000110100001011000010010000011100000101000000110000000;
        @(posedge clk) din=128'b10011111100111101001110110011100100110111001101010011001100110001001011110010110100101011001010010010011100100101001000110010000;
        @(posedge clk) din=128'b10101111101011101010110110101100101010111010101010101001101010001010011110100110101001011010010010100011101000101010000110100000;
        @(posedge clk) din=128'b10111111101111101011110110111100101110111011101010111001101110001011011110110110101101011011010010110011101100101011000110110000;
        @(posedge clk) din=128'b11001111110011101100110111001100110010111100101011001001110010001100011111000110110001011100010011000011110000101100000111000000;
        @(posedge clk) din=128'b11011111110111101101110111011100110110111101101011011001110110001101011111010110110101011101010011010011110100101101000111010000;
        @(posedge clk) din=128'b11101111111011101110110111101100111010111110101011101001111010001110011111100110111001011110010011100011111000101110000111100000;
        @(posedge clk) din=128'b11111111111111101111110111111100111110111111101011111001111110001111011111110110111101011111010011110011111100101111000111110000;

        $finish;
    end
    
    systolic_input_buffer #(
		.DATA_WIDTH(DATA_WIDTH),
		.length(length)
    ) u_systolic_input_buffer (
		.clk(clk),
		.rstn(rstn),
		.din(din),
		
		.dout(dout)
    );
    
endmodule
